module hello();
    initial 
    begin    
        $display("Hello Digital World");
    end
endmodule